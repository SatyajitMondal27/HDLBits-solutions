/*Implement the following circuit:*/
module top_module (
    output out);
supply0 gnd;
    assign out=gnd;
endmodule
