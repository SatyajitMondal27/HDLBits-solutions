/*By now, you're familiar with a module, which is a circuit that interacts with its outside through
input and output ports. Larger, more complex circuits are built by composing bigger modules out of
smaller modules and other pieces (such as assign statements and always blocks) connected together.
This forms a hierarchy, as modules can contain instances of other modules.

The figure below shows a very simple circuit with a sub-module.
 In this exercise, create one instance of module mod_a, then connect the module's three 
 pins (in1, in2, and out) to your top-level module's three ports (wires a, b, and out). 
 The module mod_a is provided for you — you must instantiate it.

When connecting modules, only the ports on the module are important. 
You do not need to know the code inside the module. 
The code for module mod_a looks like this:

Module moda.png
module mod_a ( input in1, input in2, output out );
    // Module body
endmodule
The hierarchy of modules is created by instantiating one module inside another, 
as long as all of the modules used belong to the same project (so the compiler knows where to find the module).
 The code for one module is not written inside another module's body (Code for different modules are not nested).

You may connect signals to the module by port name or port position. For extra practice, try both methods.*/
module top_module ( input a, input b, output out );
    mod_a g1(a,b,out);
endmodule
